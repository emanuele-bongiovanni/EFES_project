library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.std_logic_unsigned.all;

package mypackage is
    constant THRESHOLD_VALUE            : integer := 32;
    constant SENSING_CNT                : integer := 8;
    constant TURNING_CNT                : integer := 8;
    constant RESOLUTION                 : integer := 8;

end package mypackage;